module glib

pub type DestroyNotify fn(voidptr) voidptr
