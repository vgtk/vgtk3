module gdk
