module gtk

#pkgconfig gtk+-3.0 harfbuzz
