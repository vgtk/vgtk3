// /home/randy/code/gtk3-v/gtk3 module header

module gtk3


