module pango

pub struct Underline {
	c &PangoUnderline
}
