module gio
