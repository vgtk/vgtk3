module glib
