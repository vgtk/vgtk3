module gtk

#pkgconfig gtk+-3.0
#pkgconfig harfbuzz
