module gtk

pub struct RequestedSize {
	c &GtkRequestedSize
}
