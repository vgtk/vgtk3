module gdk

#pkgconfig gdk-3.0
#include <gdk/gdk.h>
