module gio

pub struct C.GActionGroup {}
