module gdk

pub type WindowType int

const (
	WINDOW_ROOT			= WindowType(C.GDK_WINDOW_ROOT)
	WINDOW_TOPLEVEL		= WindowType(C.GDK_WINDOW_TOPLEVEL)
	WINDOW_CHILD		= WindowType(C.GDK_WINDOW_CHILD)
	WINDOW_TEMP			= WindowType(C.GDK_WINDOW_TEMP)
	WINDOW_FOREIGN		= WindowType(C.GDK_WINDOW_FOREIGN)
	WINDOW_OFFSCREEN	= WindowType(C.GDK_WINDOW_OFFSCREEN)
	WINDOW_SUBSURFACE	= WindowType(C.GDK_WINDOW_SUBSURFACE)
)

pub type Gravity int

pub const (
	GRAVITY_NORTH_WEST = Gravity(C.GDK_GRAVITY_NORTH_WEST)
	GRAVITY_NORTH      = Gravity(C.GDK_GRAVITY_NORTH)
	GRAVITY_NORTH_EAST = Gravity(C.GDK_GRAVITY_NORTH_EAST)
	GRAVITY_WEST       = Gravity(C.GDK_GRAVITY_WEST)
	GRAVITY_CENTER     = Gravity(C.GDK_GRAVITY_CENTER)
	GRAVITY_EAST       = Gravity(C.GDK_GRAVITY_EAST)
	GRAVITY_SOUTH_WEST = Gravity(C.GDK_GRAVITY_SOUTH_WEST)
	GRAVITY_SOUTH      = Gravity(C.GDK_GRAVITY_SOUTH)
	GRAVITY_SOUTH_EAST = Gravity(C.GDK_GRAVITY_SOUTH_EAST)
	GRAVITY_STATIC     = Gravity(C.GDK_GRAVITY_STATIC)
)

pub type WindowState int

const (
	WINDOW_STATE_WITHDRAWN        = WindowState(C.GDK_WINDOW_STATE_WITHDRAWN)
	WINDOW_STATE_ICONIFIED        = WindowState(C.GDK_WINDOW_STATE_ICONIFIED)
	WINDOW_STATE_MAXIMIZED        = WindowState(C.GDK_WINDOW_STATE_MAXIMIZED)
	WINDOW_STATE_STICKY           = WindowState(C.GDK_WINDOW_STATE_STICKY)
	WINDOW_STATE_FULLSCREEN       = WindowState(C.GDK_WINDOW_STATE_FULLSCREEN)
	WINDOW_STATE_ABOVE            = WindowState(C.GDK_WINDOW_STATE_ABOVE)
	WINDOW_STATE_BELOW            = WindowState(C.GDK_WINDOW_STATE_BELOW)
	WINDOW_STATE_FOCUSED          = WindowState(C.GDK_WINDOW_STATE_FOCUSED)
	WINDOW_STATE_TILED            = WindowState(C.GDK_WINDOW_STATE_TILED)
	WINDOW_STATE_TOP_TILED        = WindowState(C.GDK_WINDOW_STATE_TOP_TILED)
	WINDOW_STATE_TOP_RESIZABLE    = WindowState(C.GDK_WINDOW_STATE_TOP_RESIZABLE)
	WINDOW_STATE_RIGHT_TILED      = WindowState(C.GDK_WINDOW_STATE_RIGHT_TILED)
	WINDOW_STATE_RIGHT_RESIZABLE  = WindowState(C.GDK_WINDOW_STATE_RIGHT_RESIZABLE)
	WINDOW_STATE_BOTTOM_TILED     = WindowState(C.GDK_WINDOW_STATE_BOTTOM_TILED)
	WINDOW_STATE_BOTTOM_RESIZABLE = WindowState(C.GDK_WINDOW_STATE_BOTTOM_RESIZABLE)
	WINDOW_STATE_LEFT_TILED       = WindowState(C.GDK_WINDOW_STATE_LEFT_TILED)
	WINDOW_STATE_LEFT_RESIZABLE   = WindowState(C.GDK_WINDOW_STATE_LEFT_RESIZABLE)
)

pub type FullScreenMode int

const (
	FULLSCREEN_ON_CURRENT_MONITOR	= FullScreenMode(C.GDK_FULLSCREEN_ON_CURRENT_MONITOR)
	FULLSCREEN_ON_ALL_MONITORS		= FullScreenMode(C.GDK_FULLSCREEN_ON_ALL_MONITORS)
)

pub type AnchorHints int

const (
	ANCHOR_FLIP_X   = AnchorHints(C.GDK_ANCHOR_FLIP_X)
	ANCHOR_FLIP_Y   = AnchorHints(C.GDK_ANCHOR_FLIP_Y)
	ANCHOR_SLIDE_X  = AnchorHints(C.GDK_ANCHOR_SLIDE_X)
	ANCHOR_SLIDE_Y  = AnchorHints(C.GDK_ANCHOR_SLIDE_Y)
	ANCHOR_RESIZE_X = AnchorHints(C.GDK_ANCHOR_RESIZE_X)
	ANCHOR_RESIZE_Y = AnchorHints(C.GDK_ANCHOR_RESIZE_Y)
	ANCHOR_FLIP     = AnchorHints(C.GDK_ANCHOR_FLIP)
	ANCHOR_SLIDE    = AnchorHints(C.GDK_ANCHOR_SLIDE)
	ANCHOR_RESIZE   = AnchorHints(C.GDK_ANCHOR_RESIZE)
)

pub type WindowEdge int

const (
	WINDOW_EDGE_NORTH_WEST = WindowEdge(C.GDK_WINDOW_EDGE_NORTH_WEST)
	WINDOW_EDGE_NORTH      = WindowEdge(C.GDK_WINDOW_EDGE_NORTH)
	WINDOW_EDGE_NORTH_EAST = WindowEdge(C.GDK_WINDOW_EDGE_NORTH_EAST)
	WINDOW_EDGE_WEST       = WindowEdge(C.GDK_WINDOW_EDGE_WEST)
	WINDOW_EDGE_EAST       = WindowEdge(C.GDK_WINDOW_EDGE_EAST)
	WINDOW_EDGE_SOUTH_WEST = WindowEdge(C.GDK_WINDOW_EDGE_SOUTH_WEST)
	WINDOW_EDGE_SOUTH      = WindowEdge(C.GDK_WINDOW_EDGE_SOUTH)
	WINDOW_EDGE_SOUTH_EAST = WindowEdge(C.GDK_WINDOW_EDGE_SOUTH_EAST)
)

pub type WindowHints int

const (
	HINT_POS         = WindowHints(C.GDK_HINT_POS)
	HINT_MIN_SIZE    = WindowHints(C.GDK_HINT_MIN_SIZE)
	HINT_MAX_SIZE    = WindowHints(C.GDK_HINT_MAX_SIZE)
	HINT_BASE_SIZE   = WindowHints(C.GDK_HINT_BASE_SIZE)
	HINT_ASPECT      = WindowHints(C.GDK_HINT_ASPECT)
	HINT_RESIZE_INC  = WindowHints(C.GDK_HINT_RESIZE_INC)
	HINT_WIN_GRAVITY = WindowHints(C.GDK_HINT_WIN_GRAVITY)
	HINT_USER_POS    = WindowHints(C.GDK_HINT_USER_POS)
	HINT_USER_SIZE   = WindowHints(C.GDK_HINT_USER_SIZE)
)

pub enum ModifierType {
	shift_mask    = 1
	lock_mask     = 2
	control_mask  = 4
	mod1_mask     = 8
	mod2_mask     = 16
	mod3_mask     = 32
	mod4_mask     = 64
	mod5_mask     = 128
	button1_mask  = 256
	button2_mask  = 512
	button3_mask  = 1024
	button4_mask  = 2048
	button5_mask  = 4096
	super_mask    = 67108864
	hyper_mask    = 134217728
	meta_mask     = 268435456
	release_mask  = 1073741824
	modifier_mask = 0x5c001fff
}

pub enum ModifierIntent {
	primary_accelerator
	context_menu
	extend_selection
	modify_selection
	no_text_input
	shift_group
	default_mod_mask
}

pub struct Window {
	c &GdkWindow
}

pub fn (w Window) get_cptr() &GdkWindow {
	return w.c
}
