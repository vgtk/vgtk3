module glib

#include <gmodule.h>
