module glib

pub type glib__CompareFn 		fn(voidptr, voidptr) int
pub type glib__CompareDataFn	fn(voidptr, voidptr, voidptr) int
