module glib

pub type CopyFunc = fn(src voidptr, data voidptr) voidptr
