module gtk

pub struct RequestedSize {
	c &C.GtkRequestedSize
}
