module pango

pub enum Style {
	normal = C.PANGO_STYLE_NORMAL
	oblique = C.PANGO_STYLE_OBLIQUE
	italic = C.PANGO_STYLE_ITALIC
}
