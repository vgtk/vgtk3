module pango

pub struct Stretch {
	c &PangoStretch
}
