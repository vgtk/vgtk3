module pango

pub struct Weight {
	c &PangoWeight
}
