module gtk

pub enum Justify {
	left
	right
	center
	fill
}

pub enum IconSize {
	invalid
	menu
	small_toolbar
	large_toolbar
	button
	dnd
	dialog
}

pub enum ReliefStyle {
	normal
	half
	@none
}
