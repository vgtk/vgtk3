module pango

pub enum Style {
	normal
	oblique
	italic
}
