module gtk

// pub struct ColorChooser {
// 	c &C.GtkColorChooser
// }

// // TODO
// pub fn (c ColorChooser) get_rgba() &C.GdkRGBA {
// 	color := &C.GdkRGBA(0)
// 	C.gtk_color_chooser_get_rgba(c.c, &color)
// 	return color
// }

// // TODO
// pub fn (c ColorChooser) set_rgba(color &C.GdkRGBA) {
// 	C.gtk_color_chooser_set_rgba(c.c, color)
// }

// pub fn (c ColorChooser) get_use_alpha() bool {
// 	return C.gtk_color_chooser_get_use_alpha(c.c)
// }

// pub fn (c ColorChooser) set_use_alpha(use_alpha bool) {
// 	C.gtk_color_chooser_set_use_alpha(c.c, use_alpha)
// }

// // TODO
// pub fn (c ColorChooser) add_palette(orientation int/* Orientation */, colors_per_line int, colors []&C.GdkRGBA) {
// 	C.gtk_color_chooser_add_palette(c.c, orientation, colors_per_line, colors.len, colors.data)
// }
