module gtk

pub enum Justify {
	left
	right
	center
	fill
}
