module gtk
#flag `pkg-config --cflags gtk+-3.0` `pkg-config --libs gtk+-3.0`
