module pango

pub struct Language {
	c &PangoLanguage
}
