module glib

pub struct C.GList
