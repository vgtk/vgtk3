module glib

pub type glib__DestroyNotify fn(voidptr) voidptr
