module gtk

pub enum ImageType {
	empty
	pixbuf
	stock
	icon_set
	animation
	icon_name
	gicon
	surface
}
