module gdk

pub type EventMask int

const (
	EXPOSURE_MASK            = EventMask(C.GDK_EXPOSURE_MASK)
	POINTER_MOTION_MASK      = EventMask(C.GDK_POINTER_MOTION_MASK)
	POINTER_MOTION_HINT_MASK = EventMask(C.GDK_POINTER_MOTION_HINT_MASK)
	BUTTON_MOTION_MASK       = EventMask(C.GDK_BUTTON_MOTION_MASK)
	BUTTON1_MOTION_MASK      = EventMask(C.GDK_BUTTON1_MOTION_MASK)
	BUTTON2_MOTION_MASK      = EventMask(C.GDK_BUTTON2_MOTION_MASK)
	BUTTON3_MOTION_MASK      = EventMask(C.GDK_BUTTON3_MOTION_MASK)
	BUTTON_PRESS_MASK        = EventMask(C.GDK_BUTTON_PRESS_MASK)
	BUTTON_RELEASE_MASK      = EventMask(C.GDK_BUTTON_RELEASE_MASK)
	KEY_PRESS_MASK           = EventMask(C.GDK_KEY_PRESS_MASK)
	KEY_RELEASE_MASK         = EventMask(C.GDK_KEY_RELEASE_MASK)
	ENTER_NOTIFY_MASK        = EventMask(C.GDK_ENTER_NOTIFY_MASK)
	LEAVE_NOTIFY_MASK        = EventMask(C.GDK_LEAVE_NOTIFY_MASK)
	FOCUS_CHANGE_MASK        = EventMask(C.GDK_FOCUS_CHANGE_MASK)
	STRUCTURE_MASK           = EventMask(C.GDK_STRUCTURE_MASK)
	PROPERTY_CHANGE_MASK     = EventMask(C.GDK_PROPERTY_CHANGE_MASK)
	VISIBILITY_NOTIFY_MASK   = EventMask(C.GDK_VISIBILITY_NOTIFY_MASK)
	PROXIMITY_IN_MASK        = EventMask(C.GDK_PROXIMITY_IN_MASK)
	PROXIMITY_OUT_MASK       = EventMask(C.GDK_PROXIMITY_OUT_MASK)
	SUBSTRUCTURE_MASK        = EventMask(C.GDK_SUBSTRUCTURE_MASK)
	SCROLL_MASK              = EventMask(C.GDK_SCROLL_MASK)
	TOUCH_MASK               = EventMask(C.GDK_TOUCH_MASK)
	SMOOTH_SCROLL_MASK       = EventMask(C.GDK_SMOOTH_SCROLL_MASK)
	TOUCHPAD_GESTURE_MASK    = EventMask(C.GDK_TOUCHPAD_GESTURE_MASK)
	TABLET_PAD_MASK          = EventMask(C.GDK_TABLET_PAD_MASK)
	ALL_EVENTS_MASK          = EventMask(C.GDK_ALL_EVENTS_MASK)
)

pub type WMDecoration int

const (
	DECOR_ALL      = WMDecoration(C.GDK_DECOR_ALL)
	DECOR_BORDER   = WMDecoration(C.GDK_DECOR_BORDER)
	DECOR_RESIZEH  = WMDecoration(C.GDK_DECOR_RESIZEH)
	DECOR_TITLE    = WMDecoration(C.GDK_DECOR_TITLE)
	DECOR_MENU     = WMDecoration(C.GDK_DECOR_MENU)
	DECOR_MINIMIZE = WMDecoration(C.GDK_DECOR_MINIMIZE)
	DECOR_MAXIMIZE = WMDecoration(C.GDK_DECOR_MAXIMIZE)
)

pub type WMFunction int

const (
	FUNC_ALL      = WMFunction(C.GDK_FUNC_ALL)
	FUNC_RESIZE   = WMFunction(C.GDK_FUNC_RESIZE)
	FUNC_MOVE     = WMFunction(C.GDK_FUNC_MOVE)
	FUNC_MINIMIZE = WMFunction(C.GDK_FUNC_MINIMIZE)
	FUNC_MAXIMIZE = WMFunction(C.GDK_FUNC_MAXIMIZE)
	FUNC_CLOSE    = WMFunction(C.GDK_FUNC_CLOSE)
)
