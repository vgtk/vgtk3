module gio

#pkgconfig gio-2.0
