module pango

pub struct FontDescription {
	c &PangoFontDescription
}
