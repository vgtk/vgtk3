module glib

pub type glib__CopyFunc fn(src voidptr, data voidptr) voidptr
