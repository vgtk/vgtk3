module glib

#pkgconfig glib-2.0
