module pango
