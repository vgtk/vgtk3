module pango

pub struct Variant {
	c &PangoVariant
}
